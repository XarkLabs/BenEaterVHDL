--
-- Based on Ben Eater's build of the SAP breadboard computer and his excellent videos.
-- https://eater.net/
--
-- Copyright (c) 2017 Ken Jordan
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.
-- 
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY counter4 IS
    PORT(
        clk_i       : IN    STD_LOGIC;
        clk_en_i    : IN    STD_LOGIC;
        rst_i       : IN    STD_LOGIC;
        set_i       : IN    STD_LOGIC;
        inc_i       : IN    STD_LOGIC;
        value_i     : IN    UNSIGNED(3 downto 0);
        value_o     : OUT   UNSIGNED(3 downto 0)
    );
END counter4;

ARCHITECTURE RTL OF counter4 IS

    SIGNAL  value   : UNSIGNED(3 downto 0) := (others => '0');

BEGIN

    PROCESS(rst_i, clk_i)
    BEGIN
        if (rst_i = '1') then
            value <= (others => '0');
        elsif (rising_edge(clk_i)) then
            if (clk_en_i = '1') then
                if (inc_i = '1') then
                    value <= value + 1;
                end if;
                if (set_i = '1') then
                    value <= value_i;
                end if;
            end if;
        end if;
    END PROCESS;
    
    value_o <= value;
    
END ARCHITECTURE RTL;
